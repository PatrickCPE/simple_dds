module wb_interface (/*AUTOARG*/
   // Outputs
   wb_dat_o, wb_ack_o, map_wr_en_o, map_wr_addr_o, map_wr_dat_o, mem_wr_en_o,
   mem_wr_addr_o, mem_wr_dat_o,
   // Inputs
   wb_clk_i, wb_rst_i, wb_dat_i, wb_addr_i, wb_lock_i, wb_cyc_i, wb_we_i
   ) ;
   //------------------------------------------------------------------------------------------------------------------------
   // Parameters
   //------------------------------------------------------------------------------------------------------------------------
   parameter DATA_WIDTH = 32;
   parameter ADDR_WIDTH = 5;
   parameter WAVE_WIDTH = 16;

   //------------------------------------------------------------------------------------------------------------------------
   // I/O
   //------------------------------------------------------------------------------------------------------------------------
   // Wishbone Interface Signals
   input wire wb_clk_i;
   input wire wb_rst_i;
   input wire [DATA_WIDTH-1:0] wb_dat_i;
   input wire [ADDR_WIDTH-1:0] wb_addr_i;
   input wire                  wb_lock_i;
   input wire                  wb_cyc_i;
   input wire                  wb_we_i;

   output wire [DATA_WIDTH-1:0] wb_dat_o;
   output wire                  wb_ack_o;


   output wire                  map_wr_en_o;
   output wire [ADDR_WIDTH-1:0] map_wr_addr_o;
   output wire [DATA_WIDTH-1:0] map_wr_dat_o;

   output wire                  mem_wr_en_o;
   output wire [ADDR_WIDTH-1:0] mem_wr_addr_o;
   output wire [DATA_WIDTH-1:0] mem_wr_dat_o;

   //------------------------------------------------------------------------------------------------------------------------
   // Internal Signals
   //------------------------------------------------------------------------------------------------------------------------

   //------------------------------------------------------------------------------------------------------------------------
   // Module Instantiations
   //------------------------------------------------------------------------------------------------------------------------

   //------------------------------------------------------------------------------------------------------------------------
   // RTL
   //------------------------------------------------------------------------------------------------------------------------
   always @ (posedge wb_clk_i) begin
      if(wb_rst_i) begin
         // TODO reset any internal registers
         wb_ack_o <= 1'b0;
      end else begin
      end
   end

   //------------------------------------------------------------------------------------------------------------------------
   // Assigns
   //------------------------------------------------------------------------------------------------------------------------

endmodule // wb_interface
